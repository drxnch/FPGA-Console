library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_ARITH.all;
use IEEE.STD_LOGIC_SIGNED.all;

entity bird is
  port (
    clk, click              : in std_logic;
    pixel_row, pixel_column : in std_logic_vector(9 downto 0);
    bird_on                 : out std_logic;
    rgb_bird                : out std_logic_vector(23 downto 0)
  );
end entity bird;

architecture behaviour of bird is

  signal size          : std_logic_vector(9 downto 0)  := conv_std_logic_vector(8, 10); -- Size of bird
  signal bird_y_pos    : std_logic_vector(9 downto 0)  := CONV_STD_LOGIC_VECTOR(240, 8);
  signal bird_x_pos    : std_logic_vector(10 downto 0) := conv_std_logic_vector(150, 11); -- x-position on of bird (compared to VGA's 640 pixels)
  signal bird_y_motion : std_logic_vector(9 downto 0)  := "0000000010";
  signal bird_x_motion : std_logic_vector(10 downto 0) := "00000000010";
  signal v_bird_on     : std_logic;
  signal u_rom_mux_out : std_logic_vector(12 downto 0); -- 1-bit alpha and 12-bit color

begin

  -- Moving bird mechanism
  Move_bird : process (click, clk)
    variable previousYbirdMotion : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR(0, 10);
    -- variable left_click_pressed  : std_logic                    := '0';
  begin
    if (rising_edge(clk)) then
      -- Apply gravity effect
      if (click = '0') then -- Check if left click is pressed
        bird_y_motion <= previousYbirdMotion + conv_std_logic_vector(1, 10); -- Increase downward motion
        if (bird_y_motion = conv_std_logic_vector(15, 10)) then
          bird_y_motion <= conv_std_logic_vector(15, 10);
        end if;

        -- Check if left click is active (jump)
      elsif (click = '1') then
        -- Apply upward impulse for a short duration
        bird_y_motion <= - CONV_STD_LOGIC_VECTOR(7, 10); -- Set initial upward motion

      end if;

      --Condition if bird hits ground
      if (('0' & bird_y_pos >= CONV_STD_LOGIC_VECTOR(450, 10) - size)) then
        bird_y_motion           <= - CONV_STD_LOGIC_VECTOR(1, 10);
      elsif ('0' & bird_y_pos <= size + 8) then
        bird_y_motion           <= CONV_STD_LOGIC_VECTOR(1, 10);
      end if;

      -- Update bird position
      bird_y_pos <= bird_y_pos + bird_y_motion;

      -- Update previous motion for next iteration
      previousYbirdMotion := bird_y_motion;
    end if;
  end process;

  SPRITE : process (v_bird_on, pixel_column, pixel_row)
    variable temp_c    : unsigned(10 downto 0) := (others => '0');
    variable temp_r    : unsigned(9 downto 0)  := (others => '0');
    variable half_size : std_logic_vector(8 downto 0);
  begin

    -- Displaying the position of bird for priority_controller to draw
    if ('0' & bird_x_pos <= '0' & pixel_column + size) and ('0' & pixel_column <= '0' & bird_x_pos + size) and
      ('0' & bird_y_pos <= pixel_row + size) and ('0' & pixel_row <= bird_y_pos + size) then
      v_bird_on <= '1';
    else
      v_bird_on <= '0';
    end if;

    half_size := size(8 downto 1) & '0';
    if (v_bird_on = '1') then
      temp_c := unsigned(pixel_column) - unsigned(bird_x_pos) - unsigned(half_size);
      temp_r := unsigned(pixel_row) - unsigned(bird_y_pos) - unsigned(half_size);
    else
      temp_c := (others => '0');
      temp_r := (others => '0');
    end if;
  end process;

  bird_on  <= v_bird_on;
  rgb_bird <= (others => '1');
end behaviour;